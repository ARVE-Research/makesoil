netcdf soildata_calculated {

dimensions:
	x = 2340 ;
	y = 2700 ;
  depth = UNLIMITED ;
  nb = 2 ;

variables:

	double x(x) ;
		x:standard_name = "projection_x_coordinate" ;
		x:units = "meter" ;
		x:axis = "X" ;
		x:actual_range = 0.,0. ;
		x:axis = "X" ;
		x:_Storage = "contiguous" ;

	double y(y) ;
		y:standard_name = "projection_y_coordinate" ;
		y:units = "meter" ;
		y:axis = "Y" ;
		y:actual_range = 0.,0. ;
		y:axis = "Y" ;
		y:_Storage = "contiguous" ;

	double lon(y, x) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:actual_range = -180., 180. ;
		lon:grid_mapping = "crs" ;

	double lat(y, x) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:actual_range = -90., 90. ;
		lat:grid_mapping = "crs" ;

  float depth(depth) ;
    depth:long_name = "vertical position of layer midpoint (below soil surface)" ;
    depth:units = "cm" ;
    depth:positive = "down" ;
    depth:bounds = "layer_bnds" ;
    depth:axis = "Z" ;
    
  float layer_bnds(depth,nb) ;
    layer_bnds:units = "cm" ;
    layer_bnds:positive = "down" ;

  float dz(depth) ;
    dz:long_name = "soil layer thickness" ;
    dz:units = "cm" ;

  byte USDA(y, x) ;
    USDA:long_name = "Predicted USDA 2014 suborder classes" ;
    USDA:units = "class" ;
    USDA:_FillValue = -1b ;
    USDA:missing_value = -1b ;
    USDA:actual_range = 0b, -1b ;
    USDA:valid_range = 1b, 99b ;
    USDA:source = "SoilGrids 2017" ;
    USDA:_Storage = "chunked" ;
    USDA:_ChunkSizes = 675, 585 ;
    USDA:_DeflateLevel = 1 ;

  short thickness(y, x) ;
    thickness:long_name = "average soil and sedimentary deposit thickness" ;
    thickness:units = "m" ;
    thickness:_FillValue = -32768s ;
    thickness:missing_value = -32768s ;
    thickness:actual_range = 100.f, -100.f ;
    thickness:scale_factor = 0.001f ;
    thickness:add_offset = 32.767f ;
    thickness:source = "Pelletier et al., 2016" ;
    thickness:_Shuffle = "true" ;
    thickness:_Storage = "chunked" ;
    thickness:_ChunkSizes = 675, 585 ;
    thickness:_DeflateLevel = 1 ;
    
  short sand(depth, y, x) ;
    sand:long_name = "sand content by mass" ;
    sand:units = "fraction" ;
    sand:_FillValue = -32768s ;
    sand:missing_value = -32768s ;
    sand:actual_range = 100.f, -100.f ;
    sand:valid_range = 0s, 1000s ;
    sand:scale_factor = 0.001f ;
    sand:source = "SoilGrids 2020" ;
    sand:_Shuffle = "true" ;
    sand:_Storage = "chunked" ;
    sand:_ChunkSizes = 1, 675, 585 ;
    sand:_DeflateLevel = 1 ;

  short clay(depth, y, x) ;
    clay:long_name = "clay content by mass" ;
    clay:units = "fraction" ;
    clay:_FillValue = -32768s ;
    clay:missing_value = -32768s ;
    clay:actual_range = 100.f, -100.f ;
    clay:valid_range = 0s, 1000s ;
    clay:scale_factor = 0.001f ;
    clay:source = "SoilGrids 2020" ;
    clay:_Shuffle = "true" ;
    clay:_Storage = "chunked" ;
    clay:_ChunkSizes = 1, 675, 585 ;
    clay:_DeflateLevel = 1 ;

  short cfvo(depth, y, x) ;
    cfvo:long_name = "coarse fragments by volume" ;
    cfvo:units = "fraction" ;
    cfvo:_FillValue = -32768s ;
    cfvo:missing_value = -32768s ;
    cfvo:actual_range = 100.f, -100.f ;
    cfvo:valid_range = 0s, 1000s ;
    cfvo:scale_factor = 0.001f ;
    cfvo:source = "SoilGrids 2020" ;
    cfvo:_Shuffle = "true" ;
    cfvo:_Storage = "chunked" ;
    cfvo:_ChunkSizes = 1, 675, 585 ;
    cfvo:_DeflateLevel = 1 ;

  short soc(depth, y, x) ;
    soc:long_name = "Soil organic carbon content by mass" ;
    soc:units = "fraction" ;
    soc:_FillValue = -32768s ;
    soc:missing_value = -32768s ;
    soc:actual_range = 100.f, -100.f ;
    soc:valid_range = 0s, 10000s ;
    soc:scale_factor = 0.0001f ;
    soc:source = "SoilGrids 2020" ;
    soc:_Shuffle = "true" ;
    soc:_Storage = "chunked" ;
    soc:_ChunkSizes = 1, 675, 585 ;
    soc:_DeflateLevel = 1 ;

  float bulk(depth, y, x) ;
    bulk:long_name = "calculated bulk density" ;
    bulk:units = "g cm-3" ;
    bulk:_FillValue = -9999.f ;
    bulk:missing_value = -9999.f ;
    bulk:actual_range = 100.f, -100.f ;
    bulk:source = "Balland et al., 2008" ;
    bulk:_Storage = "chunked" ;
    bulk:_ChunkSizes = 1, 675, 585 ;
    bulk:_DeflateLevel = 1 ;

  float Tsat(depth, y, x) ;
    Tsat:long_name = "soil porosity (Theta-sat)" ;
    Tsat:units = "fraction" ;
    Tsat:_FillValue = -9999.f ;
    Tsat:missing_value = -9999.f ;
    Tsat:actual_range = 100.f, -100.f ;
    Tsat:source = "Sandoval et al., 2024" ;
    Tsat:_Storage = "chunked" ;
    Tsat:_ChunkSizes = 1, 675, 585 ;
    Tsat:_DeflateLevel = 1 ;

  float T33(depth, y, x) ;
    T33:long_name = "soil water content at field capacity (-33 kPa)" ;
    T33:units = "mm cm-1" ;
    T33:_FillValue = -9999.f ;
    T33:missing_value = -9999.f ;
    T33:actual_range = 100.f, -100.f ;
    T33:source = "Sandoval et al., 2024" ;
    T33:_Storage = "chunked" ;
    T33:_ChunkSizes = 1, 675, 585 ;
    T33:_DeflateLevel = 1 ;

  float T1500(depth, y, x) ;
    T1500:long_name = "soil water content at permanent wilting point (-1500 kPa)" ;
    T1500:units = "mm cm-1" ;
    T1500:_FillValue = -9999.f ;
    T1500:missing_value = -9999.f ;
    T1500:actual_range = 100.f, -100.f ;
    T1500:source = "Sandoval et al., 2024" ;
    T1500:_Storage = "chunked" ;
    T1500:_ChunkSizes = 1, 675, 585 ;
    T1500:_DeflateLevel = 1 ;

  float whc(depth, y, x) ;
    whc:long_name = "water holding capacity defined as T33-T1500, reduced for coarse fragment volume" ;
    whc:units = "mm cm-1" ;
    whc:_FillValue = -9999.f ;
    whc:missing_value = -9999.f ;
    whc:actual_range = 100.f, -100.f ;
    whc:_Storage = "chunked" ;
    whc:_ChunkSizes = 1, 675, 585 ;
    whc:_DeflateLevel = 1 ;

  float Ksat(depth, y, x) ;
    Ksat:long_name = "saturated hydraulic conductivity" ;
    Ksat:units = "mm h-1" ;
    Ksat:_FillValue = -9999.f ;
    Ksat:missing_value = -9999.f ;
    Ksat:actual_range = 100.f, -100.f ;
    Ksat:source = "Sandoval et al., 2024 (code only)" ;
    Ksat:_Storage = "chunked" ;
    Ksat:_ChunkSizes = 1, 675, 585 ;

  float lambda(depth, y, x) ;
    lambda:long_name = "pore size distribution index" ;
    lambda:units = "unitless" ;
    lambda:_FillValue = -9999.f ;
    lambda:missing_value = -9999.f ;
    lambda:actual_range = 100.f, -100.f ;
    lambda:source = "Sandoval et al., after Saxton and Rawls (2006; eqn 18)" ;
    lambda:_Storage = "chunked" ;
    lambda:_ChunkSizes = 1, 675, 585 ;

  float psi_e(depth, y, x) ;
    psi_e:long_name = "tension at air entry" ;
    psi_e:units = "mm" ;
    psi_e:_FillValue = -9999.f ;
    psi_e:missing_value = -9999.f ;
    psi_e:actual_range = 100.f, -100.f ;
    psi_e:source = "Saxton and Rawls (2006; eqn 4) (converted to mm)" ;
    psi_e:_Storage = "chunked" ;
    psi_e:_ChunkSizes = 1, 675, 585 ;

// global attributes:
    :Conventions = "CF-1.11" ;
    :title = "Primary and derived soil properties" ;
    :citation1 = "Hengl, T., Mendes de Jesus, J., Heuvelink, G. B., Ruiperez Gonzalez, M., Kilibarda, M., Blagotic, A., Shangguan, W., Wright, M. N., Geng, X., Bauer-Marschallinger, B., Guevara, M. A., Vargas, R., MacMillan, R. A., Batjes, N. H., Leenaars, J. G., Ribeiro, E., Wheeler, I., Mantel, S., & Kempen, B. (2017). SoilGrids250m: Global gridded soil information based on machine learning. PLoS One, 12(2), e0169748. doi:10.1371/journal.pone.0169748" ;
    :citation2 = "Pelletier, J. D., Broxton, P. D., Hazenberg, P., Zeng, X., Troch, P. A., Niu, G. Y., Williams, Z., Brunke, M. A., & Gochis, D. (2016). A gridded global data set of soil, intact regolith, and sedimentary deposit thicknesses for regional and global land surface modeling. Journal of Advances in Modeling Earth Systems, 8(1), 41-65. doi:10.1002/2015ms000526" ;
    :citation4 = "Balland, V., Pollacco, J. A. P., & Arp, P. A. (2008). Modeling soil hydraulic properties for a wide range of soil conditions. Ecological Modelling, 219(3-4), 300-316. doi:10.1016/j.ecolmodel.2008.07.009" ;
    :citation3 = "Sandoval, D., Prentice, I. C., & Nóbrega, R. L. B. (2024). Simple process-led algorithms for simulating habitats (SPLASH v.2.0): robust calculations of water and energy fluxes. Geoscientific Model Development, 17(10), 4229-4309. doi:10.5194/gmd-17-4229-2024" ;
    :node_offset = 1 ;

}
